package axi4_lite_package;

`include "uvm_macros.svh"
import uvm_pkg::*;

`include "axi4_lite_transaction.sv"
`include "axi4_lite_monitor.sv"
`include "axi4_lite_sequencer.sv"
`include "axi4_lite_sequencer_library.sv"
`include "axi4_lite_driver.sv"
`include "axi4_lite_agent.sv"
`include "axi4_lite_scoreboard.sv"
`include "axi4_lite_environment.sv"
`include "axi4_lite_tests.sv"

endpackage: axi4_lite_package