//`ifndef DATATYPES_SV
//`define DATATYPES_SV

///*
    //Based on this: https://docs.amd.com/r/en-US/pg195-pcie-dma/Descriptors
//*/
//package descriptor;
    //typedef struct packed {
        //logic [7:0] control,
        //logic [5:0] nxt_adj, //Number of adjacent descriptors
        //logic [1:0] rsv,
        //logic [15:0] magic,
        //logic [31:0] len, //Last 4'bit are 0
        //logic [63:0] src_adr, //source address
        //logic [63:0] dst_adr, //destination address
        //logic [63:0] nxt_adr //addres of the next descriptor
    //} descriptor; //256bits
//endpackage

//`endif
